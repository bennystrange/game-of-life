magic
tech scmos
timestamp 1744959579
<< metal1 >>
rect -1453 3327 -1449 3381
rect -1453 3323 -1347 3327
rect -1153 3146 -1149 3382
rect -854 3191 -850 3381
rect -576 3349 -572 3382
rect -341 3221 -337 3383
rect -276 3349 -272 3383
rect -41 3249 -36 3382
rect 46 3297 50 3383
rect 624 3349 628 3382
rect 859 3301 863 3383
rect 946 3283 952 3381
rect 1224 3349 1228 3382
rect 1459 3271 1464 3381
rect 1524 3349 1528 3382
rect 1761 3229 1765 3382
rect 1847 3204 1851 3382
rect 2147 3159 2151 3382
rect 2746 3126 2751 3384
rect 3046 3071 3050 3382
rect 3083 3147 3282 3151
rect 3056 2847 3283 2851
rect 3189 2548 3282 2552
rect 3213 2247 3282 2251
rect -1494 2048 -1460 2052
rect 3242 1947 3281 1951
rect 3242 1346 3282 1350
rect 3240 1046 3281 1050
rect -1481 1024 -1460 1028
rect 3231 746 3282 750
rect 3200 446 3282 451
rect -1489 247 -1460 251
rect 3140 147 3282 151
rect 3109 -454 3282 -450
rect 3076 -753 3282 -749
rect -876 -1382 -872 -1347
<< m2contact >>
rect -1453 3381 -1449 3385
rect -1153 3382 -1149 3386
rect -1347 3323 -1343 3327
rect -854 3381 -850 3385
rect -576 3382 -572 3386
rect -576 3344 -572 3349
rect -341 3383 -337 3387
rect -276 3383 -272 3387
rect -276 3344 -272 3349
rect -41 3382 -36 3386
rect 46 3383 50 3387
rect 444 3386 448 3390
rect 2542 3387 2547 3392
rect 624 3382 628 3386
rect 624 3344 628 3349
rect 859 3383 863 3387
rect 859 3297 863 3301
rect 946 3381 952 3385
rect 46 3293 50 3297
rect 1224 3382 1228 3386
rect 1224 3344 1228 3349
rect 1459 3381 1464 3385
rect 946 3279 952 3283
rect 1524 3382 1528 3386
rect 1524 3344 1528 3349
rect 1761 3382 1765 3386
rect 1459 3267 1464 3271
rect -41 3245 -36 3249
rect 1761 3225 1765 3229
rect 1847 3382 1851 3386
rect -341 3217 -337 3221
rect 1847 3200 1851 3204
rect 2147 3382 2151 3386
rect -854 3187 -850 3191
rect 2147 3155 2151 3159
rect 2746 3384 2751 3388
rect -1153 3142 -1149 3146
rect 2746 3122 2751 3126
rect 3046 3382 3050 3386
rect 3079 3147 3083 3151
rect 3282 3147 3286 3151
rect 3046 3067 3050 3071
rect 3052 2847 3056 2851
rect 3283 2847 3287 2851
rect 3185 2548 3189 2552
rect 3282 2548 3286 2552
rect 3209 2247 3213 2251
rect 3282 2247 3286 2251
rect -1460 2048 -1455 2052
rect 3238 1947 3242 1951
rect 3281 1947 3285 1951
rect 3238 1346 3242 1350
rect 3282 1346 3286 1350
rect 3236 1046 3240 1050
rect 3281 1046 3285 1050
rect -1486 1024 -1481 1028
rect -1460 1024 -1455 1028
rect 3227 746 3231 750
rect 3282 746 3286 750
rect 3196 446 3200 451
rect 3282 446 3287 451
rect -1460 247 -1455 251
rect 3282 147 3286 151
rect 3105 -454 3109 -450
rect 3282 -454 3286 -450
rect 3072 -753 3076 -749
rect 3282 -753 3286 -749
rect -876 -1347 -872 -1342
rect -876 -1386 -872 -1382
rect -155 -1389 -151 -1385
rect 1644 -1389 1648 -1385
<< metal2 >>
rect -1476 3374 -1471 3382
rect -1177 3374 -1171 3387
rect -877 3374 -871 3388
rect 23 3374 29 3386
rect 444 3374 448 3386
rect 923 3374 928 3385
rect 1823 3374 1829 3385
rect 2123 3374 2129 3385
rect 2542 3374 2547 3387
rect 2723 3374 2729 3385
rect 3023 3374 3029 3385
rect -1476 3369 3266 3374
rect -1476 3129 -1471 3369
rect -1487 3123 -1471 3129
rect -1476 2829 -1471 3123
rect -1487 2823 -1471 2829
rect -1476 2529 -1471 2823
rect -1486 2523 -1471 2529
rect -1476 2229 -1471 2523
rect -1486 2223 -1471 2229
rect -1476 1877 -1471 2223
rect -1486 1871 -1471 1877
rect -1476 1329 -1471 1871
rect -1487 1323 -1471 1329
rect -1476 729 -1471 1323
rect -1486 723 -1471 729
rect -1476 429 -1471 723
rect -1486 423 -1471 429
rect -1476 77 -1471 423
rect -1487 71 -1471 77
rect -1476 -471 -1471 71
rect -1486 -477 -1471 -471
rect -1476 -771 -1471 -477
rect -1486 -777 -1471 -771
rect -1476 -1071 -1471 -777
rect -1486 -1077 -1471 -1071
rect -1476 -1365 -1471 -1077
rect -1460 3344 -576 3349
rect -572 3344 -276 3349
rect -272 3344 624 3349
rect 628 3344 1224 3349
rect 1228 3344 1524 3349
rect -1460 2052 -1455 3344
rect -1347 3071 -1343 3323
rect 729 3297 859 3301
rect 50 3293 709 3297
rect -36 3245 693 3249
rect -337 3217 597 3221
rect -850 3187 341 3191
rect -1149 3142 269 3146
rect -1347 3067 -11 3071
rect -15 2373 -11 3067
rect 265 2374 269 3142
rect 337 2373 341 3187
rect 593 2373 597 3217
rect 689 2373 693 3245
rect 705 2373 709 3293
rect 729 2373 733 3297
rect 777 3279 946 3283
rect 952 3279 953 3283
rect 777 2373 781 3279
rect 841 3267 1459 3271
rect 841 2374 845 3267
rect 873 3225 1761 3229
rect 873 2375 877 3225
rect 961 3200 1847 3204
rect 961 2373 965 3200
rect 1432 3155 2147 3159
rect 1432 2373 1436 3155
rect 1488 3126 2751 3127
rect 1488 3122 2746 3126
rect 1488 3121 2751 3122
rect 1488 2373 1492 3121
rect 1753 3067 3046 3071
rect 1753 2374 1757 3067
rect 3079 3021 3083 3147
rect 1833 3017 3083 3021
rect 3261 3129 3266 3369
rect 3261 3123 3286 3129
rect 1833 2374 1837 3017
rect -1460 1028 -1455 2048
rect 3052 1803 3056 2847
rect 3261 2829 3266 3123
rect 3261 2823 3286 2829
rect 2263 1798 3056 1803
rect 3185 1753 3189 2548
rect 3261 2529 3266 2823
rect 3261 2523 3286 2529
rect 2263 1748 3189 1753
rect 3209 1453 3213 2247
rect 3261 2229 3266 2523
rect 3261 2223 3286 2229
rect 2263 1448 3213 1453
rect 3238 1423 3242 1947
rect 2263 1418 3242 1423
rect 3261 1929 3266 2223
rect 3261 1923 3287 1929
rect 2263 1388 3242 1393
rect 3238 1350 3242 1388
rect 3261 1329 3266 1923
rect 3261 1323 3288 1329
rect -1460 251 -1455 1024
rect 3236 1023 3240 1046
rect 2263 1018 3240 1023
rect 3261 1029 3266 1323
rect 3261 1023 3288 1029
rect 2263 998 3231 1003
rect 2263 978 3200 983
rect 2263 598 3144 603
rect 2263 548 3109 553
rect 2263 488 3076 493
rect -1460 -1342 -1455 247
rect 3072 -749 3076 488
rect 3105 -450 3109 548
rect 3140 147 3144 598
rect 3196 451 3200 978
rect 3227 750 3231 998
rect 3261 729 3266 1023
rect 3261 723 3290 729
rect 3261 429 3266 723
rect 3261 423 3296 429
rect 3261 129 3266 423
rect 3261 123 3286 129
rect 3261 -471 3266 123
rect 3261 -477 3288 -471
rect 3261 -771 3266 -477
rect 3261 -777 3288 -771
rect 3261 -1071 3266 -777
rect 3261 -1077 3287 -1071
rect -1460 -1347 -876 -1342
rect 3261 -1364 3266 -1077
rect 3261 -1365 3285 -1364
rect -1476 -1370 3285 -1365
rect -1476 -1371 -1471 -1370
rect -1481 -1377 -1471 -1371
rect -1476 -1385 -1471 -1377
rect -1177 -1387 -1171 -1370
rect -577 -1386 -571 -1370
rect -155 -1385 -151 -1370
rect 23 -1385 29 -1370
rect 323 -1385 329 -1370
rect 623 -1386 629 -1370
rect 923 -1385 929 -1370
rect 1223 -1385 1229 -1370
rect 1644 -1385 1648 -1370
rect 1823 -1386 1829 -1370
rect 2123 -1385 2129 -1370
rect 2423 -1386 2429 -1370
rect 2723 -1385 2729 -1370
rect 3023 -1387 3029 -1370
rect 3278 -1378 3285 -1370
<< m3contact >>
rect 2258 1798 2263 1803
rect 2258 1748 2263 1753
rect 2258 1448 2263 1453
rect 2258 1418 2263 1423
rect 2258 1388 2263 1393
rect 2258 1018 2263 1023
rect 2258 998 2263 1003
rect 2258 978 2263 983
rect 2258 598 2263 603
rect 2258 548 2263 553
rect 2258 488 2263 493
<< metal3 >>
rect 2257 1803 2264 1804
rect 2257 1798 2258 1803
rect 2263 1798 2264 1803
rect 2257 1797 2264 1798
rect 2257 1753 2264 1754
rect 2257 1748 2258 1753
rect 2263 1748 2264 1753
rect 2257 1747 2264 1748
rect 2257 1453 2264 1454
rect 2257 1448 2258 1453
rect 2263 1448 2264 1453
rect 2257 1447 2264 1448
rect 2257 1423 2264 1424
rect 2257 1418 2258 1423
rect 2263 1418 2264 1423
rect 2257 1417 2264 1418
rect 2257 1393 2264 1394
rect 2257 1388 2258 1393
rect 2263 1388 2264 1393
rect 2257 1387 2264 1388
rect 2257 1023 2264 1024
rect 2257 1018 2258 1023
rect 2263 1018 2264 1023
rect 2257 1017 2264 1018
rect 2257 1003 2264 1004
rect 2257 998 2258 1003
rect 2263 998 2264 1003
rect 2257 997 2264 998
rect 2257 983 2264 984
rect 2257 978 2258 983
rect 2263 978 2264 983
rect 2257 977 2264 978
rect 2257 603 2264 604
rect 2257 598 2258 603
rect 2263 598 2264 603
rect 2257 597 2264 598
rect 2257 553 2264 554
rect 2257 548 2258 553
rect 2263 548 2264 553
rect 2257 547 2264 548
rect 2257 493 2264 494
rect 2257 488 2258 493
rect 2263 488 2264 493
rect 2257 487 2264 488
use PadFC  16_0
timestamp 1681001061
transform 1 0 -2500 0 1 3400
box 327 -3 1003 673
use PadFC  16_1
timestamp 1681001061
transform 0 1 3300 -1 0 4400
box 327 -3 1003 673
use PadFC  16_2
timestamp 1681001061
transform 0 -1 -1500 1 0 -2400
box 327 -3 1003 673
use PadFC  16_3
timestamp 1681001061
transform -1 0 4300 0 -1 -1400
box 327 -3 1003 673
use PadBiDir  17_0
timestamp 1711830429
transform 1 0 -1500 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_1
timestamp 1711830429
transform 1 0 -1200 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_2
timestamp 1711830429
transform 1 0 -900 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_3
timestamp 1711830429
transform 1 0 -600 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_4
timestamp 1711830429
transform 1 0 -300 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_5
timestamp 1711830429
transform 1 0 0 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_6
timestamp 1711830429
transform 1 0 600 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_7
timestamp 1711830429
transform 1 0 900 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_8
timestamp 1711830429
transform 1 0 1200 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_9
timestamp 1711830429
transform 0 -1 -1500 1 0 3100
box -36 -19 303 1000
use PadBiDir  17_10
timestamp 1711830429
transform 0 -1 -1500 1 0 2800
box -36 -19 303 1000
use PadBiDir  17_11
timestamp 1711830429
transform 0 -1 -1500 1 0 2500
box -36 -19 303 1000
use PadBiDir  17_12
timestamp 1711830429
transform 0 -1 -1500 1 0 2200
box -36 -19 303 1000
use PadBiDir  17_13
timestamp 1711830429
transform 0 -1 -1500 -1 0 1900
box -36 -19 303 1000
use PadBiDir  17_14
timestamp 1711830429
transform 0 -1 -1500 1 0 -500
box -36 -19 303 1000
use PadBiDir  17_15
timestamp 1711830429
transform 0 -1 -1500 1 0 -800
box -36 -19 303 1000
use PadBiDir  17_16
timestamp 1711830429
transform 0 -1 -1500 1 0 -1100
box -36 -19 303 1000
use PadBiDir  17_17
timestamp 1711830429
transform 0 1 3300 1 0 3100
box -36 -19 303 1000
use PadBiDir  17_18
timestamp 1711830429
transform 0 1 3300 1 0 2800
box -36 -19 303 1000
use PadBiDir  17_19
timestamp 1711830429
transform 0 1 3300 1 0 2500
box -36 -19 303 1000
use PadBiDir  17_20
timestamp 1711830429
transform 0 1 3300 1 0 2200
box -36 -19 303 1000
use PadBiDir  17_21
timestamp 1711830429
transform 0 1 3300 1 0 1900
box -36 -19 303 1000
use PadBiDir  17_22
timestamp 1711830429
transform 0 1 3300 1 0 -500
box -36 -19 303 1000
use PadBiDir  17_23
timestamp 1711830429
transform 0 1 3300 1 0 -800
box -36 -19 303 1000
use PadBiDir  17_24
timestamp 1711830429
transform 0 1 3300 1 0 -1100
box -36 -19 303 1000
use PadBiDir  17_25
timestamp 1711830429
transform 0 -1 -1500 1 0 -1400
box -36 -19 303 1000
use PadBiDir  17_26
timestamp 1711830429
transform 1 0 -1500 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_27
timestamp 1711830429
transform 1 0 -1200 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_28
timestamp 1711830429
transform 1 0 -900 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_29
timestamp 1711830429
transform 1 0 -600 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_30
timestamp 1711830429
transform 1 0 0 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_31
timestamp 1711830429
transform 1 0 300 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_32
timestamp 1711830429
transform 1 0 600 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_33
timestamp 1711830429
transform 1 0 900 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_34
timestamp 1711830429
transform 0 1 3300 1 0 -1400
box -36 -19 303 1000
use PadBiDir  17_35
timestamp 1711830429
transform 1 0 1200 0 -1 -1400
box -36 -19 303 1000
use PadVdd  18_0
timestamp 1711831643
transform 1 0 300 0 1 3400
box -3 -16 303 1000
use PadVdd  18_1
timestamp 1711831643
transform 1 0 -300 0 -1 -1400
box -3 -16 303 1000
use PadGnd  19_0
timestamp 1711831454
transform 0 -1 -1500 -1 0 2200
box -3 -11 303 1000
use PadGnd  19_1
timestamp 1711831454
transform 0 1 3300 -1 0 1900
box -3 -11 303 1000
use PadBiDir  PadBiDir_0
timestamp 1711830429
transform 1 0 1500 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_1
timestamp 1711830429
transform 1 0 1800 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_2
timestamp 1711830429
transform 1 0 2100 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_3
timestamp 1711830429
transform 1 0 2700 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_4
timestamp 1711830429
transform 1 0 3000 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_5
timestamp 1711830429
transform 1 0 1800 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_6
timestamp 1711830429
transform 1 0 2100 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_7
timestamp 1711830429
transform 1 0 2400 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_8
timestamp 1711830429
transform 1 0 2700 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_9
timestamp 1711830429
transform 1 0 3000 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_10
timestamp 1711830429
transform 0 -1 -1500 -1 0 100
box -36 -19 303 1000
use PadBiDir  PadBiDir_11
timestamp 1711830429
transform 0 -1 -1500 1 0 400
box -36 -19 303 1000
use PadBiDir  PadBiDir_12
timestamp 1711830429
transform 0 -1 -1500 1 0 700
box -36 -19 303 1000
use PadBiDir  PadBiDir_13
timestamp 1711830429
transform 0 -1 -1500 1 0 1000
box -36 -19 303 1000
use PadBiDir  PadBiDir_14
timestamp 1711830429
transform 0 -1 -1500 1 0 1300
box -36 -19 303 1000
use PadBiDir  PadBiDir_15
timestamp 1711830429
transform 0 1 3300 1 0 100
box -36 -19 303 1000
use PadBiDir  PadBiDir_16
timestamp 1711830429
transform 0 1 3300 1 0 400
box -36 -19 303 1000
use PadBiDir  PadBiDir_17
timestamp 1711830429
transform 0 1 3300 1 0 700
box -36 -19 303 1000
use PadBiDir  PadBiDir_18
timestamp 1711830429
transform 0 1 3300 1 0 1000
box -36 -19 303 1000
use PadBiDir  PadBiDir_19
timestamp 1711830429
transform 0 1 3300 1 0 1300
box -36 -19 303 1000
use PadGnd  PadGnd_0
timestamp 1711831454
transform 0 -1 -1500 -1 0 400
box -3 -11 303 1000
use PadGnd  PadGnd_1
timestamp 1711831454
transform 0 1 3300 -1 0 100
box -3 -11 303 1000
use PadVdd  PadVdd_0
timestamp 1711831643
transform 1 0 2400 0 1 3400
box -3 -16 303 1000
use PadVdd  PadVdd_1
timestamp 1711831643
transform 1 0 1500 0 -1 -1400
box -3 -16 303 1000
use TOP_SEVEN  TOP_SEVEN_0
timestamp 1744959579
transform 1 0 -465 0 1 -264
box 0 0 2728 2640
<< end >>
