magic
tech scmos
timestamp 1745093098
<< metal1 >>
rect -1366 4182 -1339 4205
rect -1059 4181 -1033 4203
rect -761 4187 -735 4209
rect -464 4195 -438 4217
rect -165 4198 -139 4220
rect 129 4204 155 4226
rect 734 4201 760 4223
rect 1030 4204 1056 4226
rect 1336 4204 1362 4226
rect 1641 4201 1667 4223
rect 1940 4201 1966 4223
rect 2231 4201 2257 4223
rect 2836 4207 2862 4229
rect 3138 4204 3164 4226
rect -1453 3327 -1449 3381
rect -1453 3323 -1347 3327
rect -2320 3209 -2264 3299
rect -1482 3146 -1292 3150
rect -2328 2901 -2272 2991
rect -1296 2941 -1292 3146
rect -1153 3146 -1149 3382
rect -854 3191 -850 3381
rect -576 3349 -572 3382
rect -341 3221 -337 3383
rect -276 3349 -272 3383
rect -41 3249 -36 3382
rect 46 3297 50 3383
rect 624 3349 628 3382
rect 2552 3386 2554 3388
rect 859 3301 863 3383
rect 946 3283 952 3381
rect 1224 3349 1228 3382
rect 1459 3271 1464 3381
rect 1524 3349 1528 3382
rect 1761 3229 1765 3382
rect 1847 3204 1851 3382
rect 2147 3159 2151 3382
rect 2746 3126 2751 3384
rect 3046 3071 3050 3382
rect 4092 3219 4127 3274
rect 3083 3147 3282 3151
rect -1296 2937 -1222 2941
rect 4093 2912 4128 2967
rect -1482 2847 -1294 2851
rect 3056 2847 3283 2851
rect -2328 2612 -2272 2702
rect 4093 2616 4128 2671
rect -1482 2546 -1329 2550
rect 3189 2548 3282 2552
rect -2331 2315 -2275 2405
rect 4093 2310 4128 2365
rect -1482 2246 -1359 2250
rect 3213 2247 3282 2251
rect -1494 2048 -1460 2052
rect 4091 2014 4126 2069
rect 3242 1947 3281 1951
rect -1482 1849 -1406 1853
rect -2335 1707 -2279 1797
rect -2331 1407 -2275 1497
rect 4093 1423 4128 1478
rect -1482 1346 -1440 1350
rect 3242 1346 3282 1350
rect -1482 1259 -1429 1263
rect -2324 1117 -2268 1207
rect 4091 1106 4126 1161
rect 3240 1046 3281 1050
rect -1481 1024 -1460 1028
rect -2324 809 -2268 899
rect 4091 816 4126 871
rect -1482 746 -1434 750
rect 3231 746 3282 750
rect -2331 520 -2275 610
rect 4093 515 4128 570
rect -1482 447 -1396 451
rect 3200 446 3282 451
rect -1489 247 -1460 251
rect -1496 242 -1492 246
rect 4093 209 4128 264
rect 3144 147 3282 151
rect -1482 49 -1345 53
rect -2326 -100 -2270 -10
rect -422 -220 -418 -217
rect -424 -222 -418 -220
rect -424 -224 -419 -222
rect -448 -249 -443 -245
rect -2308 -390 -2252 -300
rect 4091 -383 4126 -328
rect -1482 -453 -1276 -449
rect 3109 -454 3282 -450
rect -2330 -689 -2274 -599
rect 4091 -679 4126 -624
rect -1481 -753 -1148 -749
rect 3076 -753 3282 -749
rect -2323 -996 -2267 -906
rect -1247 -1049 -1243 -825
rect -1482 -1053 -1243 -1049
rect -2317 -1286 -2261 -1196
rect -1218 -1311 -1214 -870
rect -1467 -1315 -1214 -1311
rect -1467 -1349 -1463 -1315
rect -1176 -1330 -1172 -915
rect 4096 -972 4131 -917
rect -1482 -1353 -1463 -1349
rect -1453 -1334 -1172 -1330
rect -1453 -1383 -1449 -1334
rect -1154 -1382 -1150 -991
rect 3219 -1053 3281 -1049
rect -854 -1382 -850 -1117
rect -554 -1382 -550 -1182
rect 46 -1382 50 -1216
rect 324 -1382 328 -1347
rect 559 -1382 563 -1255
rect 647 -1382 651 -1302
rect 947 -1383 951 -1332
rect 1246 -1381 1250 -1332
rect 1846 -1382 1850 -1291
rect 2146 -1381 2150 -1256
rect 2446 -1381 2450 -1215
rect 2746 -1381 2750 -1179
rect 3046 -1381 3050 -1142
rect 4093 -1288 4128 -1233
rect 3100 -1354 3283 -1350
rect -1391 -2226 -1302 -2171
rect -1089 -2218 -1000 -2163
rect -786 -2226 -697 -2171
rect -487 -2218 -398 -2163
rect 104 -2236 193 -2181
rect 396 -2233 485 -2178
rect 716 -2215 805 -2160
rect 1004 -2229 1093 -2174
rect 1293 -2226 1382 -2171
rect 1898 -2218 1987 -2163
rect 2204 -2222 2293 -2167
rect 2507 -2233 2596 -2178
rect 2806 -2240 2895 -2185
rect 3114 -2233 3203 -2178
<< m2contact >>
rect -1453 3381 -1449 3385
rect -1153 3382 -1149 3386
rect -1347 3323 -1343 3327
rect -1486 3146 -1482 3150
rect -854 3381 -850 3385
rect -576 3382 -572 3386
rect -576 3344 -572 3349
rect -341 3383 -337 3387
rect -276 3383 -272 3387
rect -276 3344 -272 3349
rect -41 3382 -36 3386
rect 46 3383 50 3387
rect 444 3386 448 3390
rect 2542 3387 2547 3392
rect 624 3382 628 3386
rect 624 3344 628 3349
rect 859 3383 863 3387
rect 859 3297 863 3301
rect 946 3381 952 3385
rect 46 3293 50 3297
rect 1224 3382 1228 3386
rect 1224 3344 1228 3349
rect 1459 3381 1464 3385
rect 946 3279 952 3283
rect 1524 3382 1528 3386
rect 1524 3344 1528 3349
rect 1761 3382 1765 3386
rect 1459 3267 1464 3271
rect -41 3245 -36 3249
rect 1761 3225 1765 3229
rect 1847 3382 1851 3386
rect -341 3217 -337 3221
rect 1847 3200 1851 3204
rect 2147 3382 2151 3386
rect -854 3187 -850 3191
rect 2147 3155 2151 3159
rect 2746 3384 2751 3388
rect -1153 3142 -1149 3146
rect 2746 3122 2751 3126
rect 3046 3382 3050 3386
rect 3079 3147 3083 3151
rect 3282 3147 3286 3151
rect 3046 3067 3050 3071
rect -1222 2937 -1218 2941
rect -1486 2847 -1482 2851
rect -1294 2847 -1290 2851
rect 3052 2847 3056 2851
rect 3283 2847 3287 2851
rect -1486 2546 -1482 2550
rect -1329 2546 -1325 2550
rect 3185 2548 3189 2552
rect 3282 2548 3286 2552
rect -1486 2246 -1482 2250
rect -1359 2246 -1355 2250
rect 3209 2247 3213 2251
rect 3282 2247 3286 2251
rect -1460 2048 -1455 2052
rect 3238 1947 3242 1951
rect 3281 1947 3285 1951
rect -1486 1849 -1482 1853
rect -1406 1849 -1402 1853
rect -1486 1346 -1482 1350
rect -1440 1346 -1436 1350
rect 3238 1346 3242 1350
rect 3282 1346 3286 1350
rect -1486 1259 -1482 1263
rect -1429 1259 -1425 1263
rect 3236 1046 3240 1050
rect 3281 1046 3285 1050
rect -1486 1024 -1481 1028
rect -1460 1024 -1455 1028
rect -1486 746 -1482 750
rect -1434 746 -1430 750
rect 3227 746 3231 750
rect 3282 746 3286 750
rect -1486 447 -1482 451
rect -1396 447 -1392 451
rect 3196 446 3200 451
rect 3282 446 3287 451
rect -1460 247 -1455 251
rect 3140 147 3144 151
rect 3282 147 3286 151
rect -1486 49 -1482 53
rect -1345 49 -1341 53
rect -1486 -453 -1482 -449
rect -1276 -453 -1272 -449
rect 3105 -454 3109 -450
rect 3282 -454 3286 -450
rect -1485 -753 -1481 -749
rect -1148 -753 -1144 -749
rect 3072 -753 3076 -749
rect 3282 -753 3286 -749
rect -1247 -825 -1243 -821
rect -1486 -1053 -1482 -1049
rect -1218 -870 -1214 -866
rect -1176 -915 -1172 -911
rect -1486 -1353 -1482 -1349
rect -1154 -991 -1150 -987
rect -1453 -1387 -1449 -1383
rect 3215 -1053 3219 -1049
rect 3281 -1053 3285 -1049
rect -1154 -1386 -1150 -1382
rect -854 -1117 -850 -1113
rect 3046 -1142 3050 -1138
rect -854 -1386 -850 -1382
rect -554 -1182 -550 -1178
rect 2746 -1179 2750 -1175
rect -554 -1386 -550 -1382
rect 46 -1216 50 -1212
rect 2446 -1215 2450 -1211
rect 559 -1255 563 -1251
rect -155 -1389 -151 -1385
rect 46 -1386 50 -1382
rect 324 -1347 328 -1342
rect 324 -1386 328 -1382
rect 2146 -1256 2150 -1252
rect 1846 -1291 1850 -1287
rect 559 -1386 563 -1382
rect 647 -1302 651 -1298
rect 647 -1386 651 -1382
rect 947 -1332 951 -1328
rect 947 -1387 951 -1383
rect 1246 -1332 1250 -1328
rect 1246 -1385 1250 -1381
rect 1644 -1389 1648 -1385
rect 1846 -1386 1850 -1382
rect 2146 -1385 2150 -1381
rect 2446 -1385 2450 -1381
rect 2746 -1385 2750 -1381
rect 3096 -1354 3100 -1350
rect 3283 -1354 3287 -1350
rect 3046 -1385 3050 -1381
<< metal2 >>
rect -1476 3374 -1471 3382
rect -1177 3374 -1171 3387
rect -877 3374 -871 3388
rect 23 3374 29 3386
rect 444 3374 448 3386
rect 923 3374 928 3385
rect 1823 3374 1829 3385
rect 2123 3374 2129 3385
rect 2542 3374 2547 3387
rect 2723 3374 2729 3385
rect 3023 3374 3029 3385
rect -1476 3369 3266 3374
rect -1476 3129 -1471 3369
rect -1487 3123 -1471 3129
rect -1476 2829 -1471 3123
rect -1487 2823 -1471 2829
rect -1476 2529 -1471 2823
rect -1486 2523 -1471 2529
rect -1476 2229 -1471 2523
rect -1486 2223 -1471 2229
rect -1476 1877 -1471 2223
rect -1486 1871 -1471 1877
rect -1476 1329 -1471 1871
rect -1487 1323 -1471 1329
rect -1476 729 -1471 1323
rect -1486 723 -1471 729
rect -1476 429 -1471 723
rect -1486 423 -1471 429
rect -1476 77 -1471 423
rect -1487 71 -1471 77
rect -1476 -471 -1471 71
rect -1486 -477 -1471 -471
rect -1476 -771 -1471 -477
rect -1486 -777 -1471 -771
rect -1476 -1071 -1471 -777
rect -1486 -1077 -1471 -1071
rect -1476 -1365 -1471 -1077
rect -1460 3344 -576 3349
rect -572 3344 -276 3349
rect -272 3344 624 3349
rect 628 3344 1224 3349
rect 1228 3344 1524 3349
rect -1460 2052 -1455 3344
rect -1347 3071 -1343 3323
rect 729 3297 859 3301
rect 50 3293 709 3297
rect -36 3245 693 3249
rect -337 3217 597 3221
rect -850 3187 341 3191
rect -1149 3142 269 3146
rect -1347 3067 -11 3071
rect -1460 1028 -1455 2048
rect -1406 1352 -1402 1849
rect -1359 1443 -1355 2246
rect -1329 1703 -1325 2546
rect -1294 1722 -1290 2847
rect -1222 1943 -1218 2937
rect -15 2373 -11 3067
rect 265 2374 269 3142
rect 337 2373 341 3187
rect 593 2373 597 3217
rect 689 2373 693 3245
rect 705 2373 709 3293
rect 729 2373 733 3297
rect 777 3279 946 3283
rect 952 3279 953 3283
rect 777 2373 781 3279
rect 841 3267 1459 3271
rect 841 2374 845 3267
rect 873 3225 1761 3229
rect 873 2375 877 3225
rect 961 3200 1847 3204
rect 961 2373 965 3200
rect 1432 3155 2147 3159
rect 1432 2373 1436 3155
rect 1488 3126 2751 3127
rect 1488 3122 2746 3126
rect 1488 3121 2751 3122
rect 1488 2373 1492 3121
rect 1753 3067 3046 3071
rect 1753 2374 1757 3067
rect 3079 3021 3083 3147
rect 1833 3017 3083 3021
rect 3261 3129 3266 3369
rect 3261 3123 3286 3129
rect 1833 2374 1837 3017
rect -1222 1939 -465 1943
rect 3052 1803 3056 2847
rect 3261 2829 3266 3123
rect 3261 2823 3286 2829
rect 2263 1798 3056 1803
rect 3185 1753 3189 2548
rect 3261 2529 3266 2823
rect 3261 2523 3286 2529
rect 2263 1748 3189 1753
rect -1294 1718 -465 1722
rect -1329 1699 -465 1703
rect 3209 1453 3213 2247
rect 3261 2229 3266 2523
rect 3261 2223 3286 2229
rect 2263 1448 3213 1453
rect -1359 1439 -465 1443
rect 3238 1423 3242 1947
rect 2263 1418 3242 1423
rect 3261 1929 3266 2223
rect 3261 1923 3287 1929
rect 2263 1388 3242 1393
rect -1406 1348 -465 1352
rect 3238 1350 3242 1388
rect -1440 1332 -1436 1346
rect -1440 1328 -465 1332
rect 3261 1329 3266 1923
rect 3261 1323 3288 1329
rect -1429 1083 -1425 1259
rect -1429 1078 -465 1083
rect -1460 251 -1455 1024
rect 3236 1023 3240 1046
rect 2263 1018 3240 1023
rect 3261 1029 3266 1323
rect 3261 1023 3288 1029
rect 2263 998 3231 1003
rect 2263 978 3200 983
rect -1434 938 -465 943
rect -1434 750 -1430 938
rect -1396 919 -465 923
rect -1396 451 -1392 919
rect -1345 869 -465 873
rect -1460 -1342 -1455 247
rect -1345 53 -1341 869
rect 2263 598 3144 603
rect 2263 548 3109 553
rect 2263 488 3076 493
rect -1276 479 -465 483
rect -1276 -449 -1272 479
rect -1148 388 -465 392
rect -1148 -749 -1144 388
rect -63 -821 -59 -264
rect -1243 -825 -59 -821
rect 25 -866 29 -264
rect -1214 -870 29 -866
rect 65 -911 69 -264
rect -1172 -915 69 -911
rect 241 -987 245 -264
rect -1150 -991 245 -987
rect 481 -1113 485 -264
rect -850 -1117 485 -1113
rect 529 -1178 533 -264
rect -550 -1182 533 -1178
rect 545 -1212 549 -264
rect 50 -1216 549 -1212
rect 913 -1251 917 -264
rect 563 -1255 917 -1251
rect 1009 -1298 1013 -264
rect 651 -1302 1013 -1298
rect 1025 -1328 1029 -264
rect 951 -1332 1029 -1328
rect 1064 -1328 1068 -264
rect 1177 -1287 1181 -264
rect 1473 -1252 1477 -264
rect 1505 -1211 1509 -264
rect 1561 -1175 1565 -264
rect 1705 -1138 1709 -264
rect 1737 -1088 1741 -264
rect 1793 -1062 1797 -264
rect 3072 -749 3076 488
rect 3105 -450 3109 548
rect 3140 151 3144 598
rect 3196 451 3200 978
rect 3227 750 3231 998
rect 3261 729 3266 1023
rect 3261 723 3290 729
rect 3261 429 3266 723
rect 3261 423 3296 429
rect 3261 129 3266 423
rect 3261 123 3286 129
rect 3261 -471 3266 123
rect 3261 -477 3288 -471
rect 3261 -771 3266 -477
rect 3261 -777 3288 -771
rect 3215 -1062 3219 -1053
rect 1793 -1066 3219 -1062
rect 3261 -1071 3266 -777
rect 3261 -1077 3287 -1071
rect 1737 -1092 3100 -1088
rect 1705 -1142 3046 -1138
rect 1561 -1179 2746 -1175
rect 1505 -1215 2446 -1211
rect 1473 -1256 2146 -1252
rect 1177 -1291 1846 -1287
rect 1064 -1332 1246 -1328
rect -1460 -1347 324 -1342
rect 3096 -1350 3100 -1092
rect 3261 -1364 3266 -1077
rect 3261 -1365 3285 -1364
rect -1476 -1370 3285 -1365
rect -1476 -1371 -1471 -1370
rect -1481 -1377 -1471 -1371
rect -1476 -1385 -1471 -1377
rect -1177 -1387 -1171 -1370
rect -876 -1386 -872 -1370
rect -577 -1386 -571 -1370
rect -155 -1385 -151 -1370
rect 23 -1385 29 -1370
rect 623 -1381 629 -1370
rect 923 -1385 929 -1370
rect 1223 -1385 1229 -1370
rect 1644 -1385 1648 -1370
rect 1823 -1386 1829 -1370
rect 2123 -1385 2129 -1370
rect 2423 -1386 2429 -1370
rect 2723 -1385 2729 -1370
rect 3023 -1387 3029 -1370
rect 3278 -1378 3285 -1370
<< m3contact >>
rect -465 1938 -460 1943
rect 2258 1798 2263 1803
rect 2258 1748 2263 1753
rect -465 1718 -460 1723
rect -465 1698 -460 1703
rect 2258 1448 2263 1453
rect -465 1438 -460 1443
rect 2258 1418 2263 1423
rect 2258 1388 2263 1393
rect -465 1348 -460 1353
rect -465 1328 -460 1333
rect -465 1078 -460 1083
rect 2258 1018 2263 1023
rect 2258 998 2263 1003
rect 2258 978 2263 983
rect -465 938 -460 943
rect -465 918 -460 923
rect -465 868 -460 873
rect 2258 598 2263 603
rect 2258 548 2263 553
rect 2258 488 2263 493
rect -465 478 -460 483
rect -465 388 -460 393
<< metal3 >>
rect -466 1943 -459 1944
rect -466 1938 -465 1943
rect -460 1938 -459 1943
rect -466 1937 -459 1938
rect 2257 1803 2264 1804
rect 2257 1798 2258 1803
rect 2263 1798 2264 1803
rect 2257 1797 2264 1798
rect 2257 1753 2264 1754
rect 2257 1748 2258 1753
rect 2263 1748 2264 1753
rect 2257 1747 2264 1748
rect -466 1723 -459 1724
rect -466 1718 -465 1723
rect -460 1718 -459 1723
rect -466 1717 -459 1718
rect -466 1703 -459 1704
rect -466 1698 -465 1703
rect -460 1698 -459 1703
rect -466 1697 -459 1698
rect 2257 1453 2264 1454
rect 2257 1448 2258 1453
rect 2263 1448 2264 1453
rect 2257 1447 2264 1448
rect -466 1443 -459 1444
rect -466 1438 -465 1443
rect -460 1438 -459 1443
rect -466 1437 -459 1438
rect 2257 1423 2264 1424
rect 2257 1418 2258 1423
rect 2263 1418 2264 1423
rect 2257 1417 2264 1418
rect 2257 1393 2264 1394
rect 2257 1388 2258 1393
rect 2263 1388 2264 1393
rect 2257 1387 2264 1388
rect -466 1353 -459 1354
rect -466 1348 -465 1353
rect -460 1348 -459 1353
rect -466 1347 -459 1348
rect -466 1333 -459 1334
rect -466 1328 -465 1333
rect -460 1328 -459 1333
rect -466 1327 -459 1328
rect -466 1083 -459 1084
rect -466 1078 -465 1083
rect -460 1078 -459 1083
rect -466 1077 -459 1078
rect 2257 1023 2264 1024
rect 2257 1018 2258 1023
rect 2263 1018 2264 1023
rect 2257 1017 2264 1018
rect 2257 1003 2264 1004
rect 2257 998 2258 1003
rect 2263 998 2264 1003
rect 2257 997 2264 998
rect 2257 983 2264 984
rect 2257 978 2258 983
rect 2263 978 2264 983
rect 2257 977 2264 978
rect -466 943 -459 944
rect -466 938 -465 943
rect -460 938 -459 943
rect -466 937 -459 938
rect -466 923 -459 924
rect -466 918 -465 923
rect -460 918 -459 923
rect -466 917 -459 918
rect -466 873 -459 874
rect -466 868 -465 873
rect -460 868 -459 873
rect -466 867 -459 868
rect 2257 603 2264 604
rect 2257 598 2258 603
rect 2263 598 2264 603
rect 2257 597 2264 598
rect 2257 553 2264 554
rect 2257 548 2258 553
rect 2263 548 2264 553
rect 2257 547 2264 548
rect 2257 493 2264 494
rect 2257 488 2258 493
rect 2263 488 2264 493
rect 2257 487 2264 488
rect -466 483 -459 484
rect -466 478 -465 483
rect -460 478 -459 483
rect -466 477 -459 478
rect -466 393 -459 394
rect -466 388 -465 393
rect -460 388 -459 393
rect -466 387 -459 388
use PadFC  16_0
timestamp 1681001061
transform 1 0 -2500 0 1 3400
box 327 -3 1003 673
use PadFC  16_1
timestamp 1681001061
transform 0 1 3300 -1 0 4400
box 327 -3 1003 673
use PadFC  16_2
timestamp 1681001061
transform 0 -1 -1500 1 0 -2400
box 327 -3 1003 673
use PadFC  16_3
timestamp 1681001061
transform -1 0 4300 0 -1 -1400
box 327 -3 1003 673
use PadBiDir  17_0
timestamp 1711830429
transform 1 0 -1500 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_1
timestamp 1711830429
transform 1 0 -1200 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_2
timestamp 1711830429
transform 1 0 -900 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_3
timestamp 1711830429
transform 1 0 -600 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_4
timestamp 1711830429
transform 1 0 -300 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_5
timestamp 1711830429
transform 1 0 0 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_6
timestamp 1711830429
transform 1 0 600 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_7
timestamp 1711830429
transform 1 0 900 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_8
timestamp 1711830429
transform 1 0 1200 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_9
timestamp 1711830429
transform 0 -1 -1500 1 0 3100
box -36 -19 303 1000
use PadBiDir  17_10
timestamp 1711830429
transform 0 -1 -1500 1 0 2800
box -36 -19 303 1000
use PadBiDir  17_11
timestamp 1711830429
transform 0 -1 -1500 1 0 2500
box -36 -19 303 1000
use PadBiDir  17_12
timestamp 1711830429
transform 0 -1 -1500 1 0 2200
box -36 -19 303 1000
use PadBiDir  17_13
timestamp 1711830429
transform 0 -1 -1500 -1 0 1900
box -36 -19 303 1000
use PadBiDir  17_14
timestamp 1711830429
transform 0 -1 -1500 1 0 -500
box -36 -19 303 1000
use PadBiDir  17_15
timestamp 1711830429
transform 0 -1 -1500 1 0 -800
box -36 -19 303 1000
use PadBiDir  17_16
timestamp 1711830429
transform 0 -1 -1500 1 0 -1100
box -36 -19 303 1000
use PadBiDir  17_17
timestamp 1711830429
transform 0 1 3300 1 0 3100
box -36 -19 303 1000
use PadBiDir  17_18
timestamp 1711830429
transform 0 1 3300 1 0 2800
box -36 -19 303 1000
use PadBiDir  17_19
timestamp 1711830429
transform 0 1 3300 1 0 2500
box -36 -19 303 1000
use PadBiDir  17_20
timestamp 1711830429
transform 0 1 3300 1 0 2200
box -36 -19 303 1000
use PadBiDir  17_21
timestamp 1711830429
transform 0 1 3300 1 0 1900
box -36 -19 303 1000
use PadBiDir  17_22
timestamp 1711830429
transform 0 1 3300 1 0 -500
box -36 -19 303 1000
use PadBiDir  17_23
timestamp 1711830429
transform 0 1 3300 1 0 -800
box -36 -19 303 1000
use PadBiDir  17_24
timestamp 1711830429
transform 0 1 3300 1 0 -1100
box -36 -19 303 1000
use PadBiDir  17_25
timestamp 1711830429
transform 0 -1 -1500 1 0 -1400
box -36 -19 303 1000
use PadBiDir  17_26
timestamp 1711830429
transform 1 0 -1500 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_27
timestamp 1711830429
transform 1 0 -1200 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_28
timestamp 1711830429
transform 1 0 -900 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_29
timestamp 1711830429
transform 1 0 -600 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_30
timestamp 1711830429
transform 1 0 0 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_31
timestamp 1711830429
transform 1 0 300 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_32
timestamp 1711830429
transform 1 0 600 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_33
timestamp 1711830429
transform 1 0 900 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_34
timestamp 1711830429
transform 0 1 3300 1 0 -1400
box -36 -19 303 1000
use PadBiDir  17_35
timestamp 1711830429
transform 1 0 1200 0 -1 -1400
box -36 -19 303 1000
use PadVdd  18_0
timestamp 1711831643
transform 1 0 300 0 1 3400
box -3 -16 303 1000
use PadVdd  18_1
timestamp 1711831643
transform 1 0 -300 0 -1 -1400
box -3 -16 303 1000
use PadGnd  19_0
timestamp 1711831454
transform 0 -1 -1500 -1 0 2200
box -3 -11 303 1000
use PadGnd  19_1
timestamp 1711831454
transform 0 1 3300 -1 0 1900
box -3 -11 303 1000
use PadBiDir  PadBiDir_0
timestamp 1711830429
transform 1 0 1500 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_1
timestamp 1711830429
transform 1 0 1800 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_2
timestamp 1711830429
transform 1 0 2100 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_3
timestamp 1711830429
transform 1 0 2700 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_4
timestamp 1711830429
transform 1 0 3000 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_5
timestamp 1711830429
transform 1 0 1800 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_6
timestamp 1711830429
transform 1 0 2100 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_7
timestamp 1711830429
transform 1 0 2400 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_8
timestamp 1711830429
transform 1 0 2700 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_9
timestamp 1711830429
transform 1 0 3000 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_10
timestamp 1711830429
transform 0 -1 -1500 -1 0 100
box -36 -19 303 1000
use PadBiDir  PadBiDir_11
timestamp 1711830429
transform 0 -1 -1500 1 0 400
box -36 -19 303 1000
use PadBiDir  PadBiDir_12
timestamp 1711830429
transform 0 -1 -1500 1 0 700
box -36 -19 303 1000
use PadBiDir  PadBiDir_13
timestamp 1711830429
transform 0 -1 -1500 1 0 1000
box -36 -19 303 1000
use PadBiDir  PadBiDir_14
timestamp 1711830429
transform 0 -1 -1500 1 0 1300
box -36 -19 303 1000
use PadBiDir  PadBiDir_15
timestamp 1711830429
transform 0 1 3300 1 0 100
box -36 -19 303 1000
use PadBiDir  PadBiDir_16
timestamp 1711830429
transform 0 1 3300 1 0 400
box -36 -19 303 1000
use PadBiDir  PadBiDir_17
timestamp 1711830429
transform 0 1 3300 1 0 700
box -36 -19 303 1000
use PadBiDir  PadBiDir_18
timestamp 1711830429
transform 0 1 3300 1 0 1000
box -36 -19 303 1000
use PadBiDir  PadBiDir_19
timestamp 1711830429
transform 0 1 3300 1 0 1300
box -36 -19 303 1000
use PadGnd  PadGnd_0
timestamp 1711831454
transform 0 -1 -1500 -1 0 400
box -3 -11 303 1000
use PadGnd  PadGnd_1
timestamp 1711831454
transform 0 1 3300 -1 0 100
box -3 -11 303 1000
use PadVdd  PadVdd_0
timestamp 1711831643
transform 1 0 2400 0 1 3400
box -3 -16 303 1000
use PadVdd  PadVdd_1
timestamp 1711831643
transform 1 0 1500 0 -1 -1400
box -3 -16 303 1000
use TOP_SEVEN  TOP_SEVEN_0
timestamp 1744959579
transform 1 0 -465 0 1 -264
box 0 0 2728 2640
<< labels >>
rlabel metal1 -1351 4192 -1351 4192 1 grid43
rlabel metal1 -1046 4191 -1046 4191 1 grid37
rlabel metal1 -749 4197 -749 4197 1 grid44
rlabel metal1 -449 4206 -449 4206 1 clkb
rlabel metal1 -150 4209 -150 4209 1 prgm
rlabel metal1 143 4211 143 4211 1 grid38
rlabel metal1 748 4210 748 4210 1 pp
rlabel metal1 1044 4214 1044 4215 1 grid45
rlabel metal1 1350 4215 1350 4215 1 btn1
rlabel metal1 1655 4212 1655 4212 1 btn0
rlabel metal1 1953 4214 1953 4214 1 grid31
rlabel metal1 2244 4209 2244 4209 1 grid46
rlabel metal1 2849 4217 2849 4217 1 grid39
rlabel metal1 3149 4212 3149 4212 1 grid47
rlabel metal1 4104 3246 4104 3246 1 grid48
rlabel metal1 4109 2940 4109 2940 1 grid40
rlabel metal1 4110 2639 4110 2639 1 grid41
rlabel metal1 4111 2340 4111 2340 1 grid32
rlabel metal1 4106 2038 4106 2038 1 grid34
rlabel metal1 4110 1450 4110 1450 1 grid33
rlabel metal1 4104 1130 4104 1130 1 grid25
rlabel metal1 4105 841 4105 841 1 grid26
rlabel metal1 4104 539 4104 539 1 grid27
rlabel metal1 4108 234 4108 234 1 grid18
rlabel metal1 4108 -359 4108 -359 1 grid20
rlabel metal1 4110 -652 4110 -652 1 grid19
rlabel metal1 4113 -947 4113 -947 1 grid12
rlabel metal1 4108 -1264 4108 -1264 1 grid13
rlabel metal1 3158 -2208 3158 -2208 1 grid5
rlabel metal1 2852 -2218 2852 -2218 1 grid6
rlabel metal1 2549 -2204 2549 -2204 1 grid11
rlabel metal1 2250 -2204 2250 -2204 1 grid4
rlabel metal1 1944 -2194 1944 -2194 1 grid3
rlabel metal1 1353 -2201 1353 -2201 1 grid10
rlabel metal1 1054 -2208 1054 -2208 1 grid24
rlabel metal1 752 -2190 752 -2190 1 grid17
rlabel metal1 445 -2208 445 -2208 1 clka
rlabel metal1 146 -2211 146 -2211 1 grid9
rlabel metal1 -437 -2190 -437 -2190 1 grid2
rlabel metal1 -740 -2204 -740 -2204 1 grid16
rlabel metal1 -1046 -2197 -1046 -2197 1 grid1
rlabel metal1 -1352 -2211 -1352 -2211 1 grid8
rlabel metal1 -2296 -1238 -2296 -1238 1 grid0
rlabel metal1 -2294 -957 -2294 -957 1 grid7
rlabel metal1 -2307 -636 -2307 -636 1 grid14
rlabel metal1 -2283 -345 -2283 -345 1 grid15
rlabel metal1 -2300 -57 -2300 -57 1 grid21
rlabel metal1 -2304 562 -2304 562 1 grid22
rlabel metal1 -2298 859 -2298 859 1 grid23
rlabel metal1 -2296 1159 -2296 1159 1 stop
rlabel metal1 -2304 1449 -2304 1449 1 grid28
rlabel metal1 -2304 1757 -2304 1757 1 grid29
rlabel metal1 -2303 2358 -2303 2358 1 grid30
rlabel metal1 -2299 2660 -2299 2660 1 grid36
rlabel metal1 -2300 2945 -2300 2945 1 grid35
rlabel metal1 -2293 3264 -2293 3264 1 grid42
rlabel metal1 2553 3387 2553 3387 1 Vdd!
rlabel metal1 -445 -247 -445 -247 1 Vdd!
rlabel metal1 -1494 244 -1494 244 1 GND!
rlabel metal1 -420 -219 -420 -219 1 GND!
<< end >>
